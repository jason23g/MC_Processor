-------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-------------------------------------------------------------------------------
ENTITY MUX_32x32_TB IS
END MUX_32x32_TB;
-------------------------------------------------------------------------------
ARCHITECTURE behavior OF MUX_32x32_TB IS

	-- Component Declaration for the Unit Under Test (UUT)
	COMPONENT MUX_32x32
	PORT (
		ctrl : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		Din0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din4 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din6 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din7 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din8 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din9 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din10 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din11 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din12 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din13 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din14 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din15 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din16 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din17 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din18 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din19 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din20 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din21 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din22 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din23 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din24 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din25 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din26 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din27 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din28 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din29 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din30 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Din31 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Dout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
	END COMPONENT; 

	--Inputs
	SIGNAL ctrl : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din0 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din1 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din2 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din3 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din4 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din5 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din6 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din7 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din8 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din9 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din10 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din11 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din12 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din13 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din14 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din15 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din16 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din17 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din18 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din19 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din20 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din21 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din22 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din23 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din24 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din25 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din26 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din27 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din28 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din29 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din30 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	SIGNAL Din31 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');

	--Outputs
	SIGNAL Dout : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	-- Instantiate the Unit Under Test (UUT)
	uut : MUX_32x32
	PORT MAP (
		ctrl => ctrl,
		Din0 => Din0,
		Din1 => Din1,
		Din2 => Din2,
		Din3 => Din3,
		Din4 => Din4,
		Din5 => Din5,
		Din6 => Din6,
		Din7 => Din7,
		Din8 => Din8,
		Din9 => Din9,
		Din10 => Din10,
		Din11 => Din11,
		Din12 => Din12,
		Din13 => Din13,
		Din14 => Din14,
		Din15 => Din15,
		Din16 => Din16,
		Din17 => Din17,
		Din18 => Din18,
		Din19 => Din19,
		Din20 => Din20,
		Din21 => Din21,
		Din22 => Din22,
		Din23 => Din23,
		Din24 => Din24,
		Din25 => Din25,
		Din26 => Din26,
		Din27 => Din27,
		Din28 => Din28,
		Din29 => Din29,
		Din30 => Din30,
		Din31 => Din31,
		Dout => Dout
	);
	
	-- Stimulus process
	stim_proc : PROCESS
	BEGIN
		-- insert stimulus here
		ctrl <= "00000";
		Din0 <= "11111111111111111100001111111111";
		WAIT FOR 100 ns;
		
		ctrl <= "00001";
		Din1 <= "11101111111000111100001111111111";
		WAIT FOR 100 ns;
		
		ctrl <= "00010";
		Din2 <= "11111000001111111100001111111111";
		WAIT FOR 100 ns;
		
		ctrl <= "00100";
		Din4 <= "11111011111111111100001111100011";
		WAIT FOR 100 ns;
		
		ctrl <= "01000";
		Din8 <= "11111111000111011100001111111111";
		WAIT FOR 100 ns;
		
		ctrl <= "10000";
		Din16 <= "00011110011111111100001111111111";
		WAIT FOR 100 ns;
		
		ctrl <= "10010";
		Din18 <= "10001111110001111000001111111101";
		WAIT FOR 100 ns;
		
		ctrl <= "11111";
		Din31 <= "10000111110011011100001111001111";
		WAIT FOR 100 ns;
		
		WAIT;
	END PROCESS;

END;
-------------------------------------------------------------------------------